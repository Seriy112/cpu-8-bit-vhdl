-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : s
-- Author      : Microsoft
-- Company     : Microsoft
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\s\s\compile\memory.vhd
-- Generated   : Fri May 13 01:12:58 2016
-- From        : c:\My_Designs\s\s\src\memory.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library ieee;
        use ieee.std_logic_1164.all;
        use ieee.std_logic_signed.all;

entity memory is
  port(
       RD : in std_logic;
       Adr : in std_logic_vector(5 downto 0);
       MrOut : out std_logic;
       InstrCom : out std_logic_vector(0 to 27)
  );
end memory;

architecture Memory of memory is

---- Architecture declarations -----
--Added by Active-HDL. Do not change code inside this section.
type MemoryType is array (0 to 59) of std_logic_vector(0 to 27);
--End of extra code.


---- Signal declarations used on the diagram ----

signal Memory : MemoryType;

begin

---- Processes ----

process (RD)
                       begin
                         if RD = '1' and RD'event then
                            InstrCom <= Memory(CONV_INTEGER('0' & Adr));
                            MrOut <= '1';
                         end if;
                         if RD = '0' and RD'event then
                            MrOut <= '0';
                         end if;
                       end process;                      

---- User Signal Assignments ----
Memory(0) <= "000" & "000000" & "0000000" & "0000000" & "0000" & "0";
Memory(1) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(2) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(3) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(4) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(5) <= "000" & "000000" & "0010000" & "0000000" & "0000" & "0";
Memory(6) <= "100" & "000000" & "0000000" & "0000000" & "0000" & "0";
Memory(7) <= "000" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(8) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(9) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(10) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(11) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(12) <= "000" & "000000" & "0000000" & "0000001" & "0000" & "0";
Memory(13) <= "001" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(14) <= "000" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(15) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(16) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(17) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(18) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(19) <= "000" & "000000" & "0000000" & "0000000" & "0010" & "0";
Memory(20) <= "000" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(21) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(22) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(23) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(24) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(25) <= "000" & "000000" & "0000000" & "0000000" & "1000" & "0";
Memory(26) <= "001" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(27) <= "000" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(28) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(29) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(30) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(31) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(32) <= "000" & "000000" & "0000000" & "0000000" & "0010" & "0";
Memory(33) <= "000" & "000000" & "0000000" & "0000000" & "0100" & "0";
Memory(34) <= "000" & "000000" & "0000000" & "0000000" & "0001" & "0";
Memory(35) <= "000" & "000000" & "0000000" & "0001000" & "0000" & "0";
Memory(36) <= "000" & "000000" & "0000000" & "0000100" & "0000" & "0";
Memory(37) <= "000" & "000000" & "0000000" & "0000001" & "0000" & "0";
Memory(38) <= "001" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(51) <= "010" & "110110" & "0000000" & "0000000" & "0000" & "0";
Memory(52) <= "000" & "000000" & "0000000" & "0000000" & "0000" & "0";
Memory(53) <= "000" & "000000" & "0000000" & "0000000" & "0000" & "0";
Memory(54) <= "000" & "000000" & "0100000" & "0000000" & "0000" & "0";
Memory(55) <= "000" & "000000" & "0001000" & "0000000" & "0000" & "0";
Memory(56) <= "000" & "000000" & "0000110" & "0000000" & "0000" & "0";
Memory(57) <= "000" & "000000" & "0000001" & "0000000" & "0000" & "0";
Memory(58) <= "000" & "000000" & "0000000" & "1000000" & "0000" & "0";
Memory(59) <= "001" & "000000" & "1000000" & "0000000" & "0000" & "0";

end Memory;
